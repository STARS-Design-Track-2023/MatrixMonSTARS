//this would be enabled from the top
