module 

endmodule